module SFT(Y,A,B,Op);
	input  [31:0] A,B;
	input  [1:0] Op;
	output [31:0] Y;

	wire [31:0]  Y1,Y2,Y3;

	LSFT  LSHIFTER  (Y1,A,B);
	RSFT  RSHIFTER  (Y2,A,B);
	ARSFT ARSHIFTER	(Y3,A,B);

assign Y= (Op==2'b00)?Y1:((Op==2'b01)?Y2:Y3);

endmodule

module LSFT(Y,A,B);
	input  [31:0] A,B;
	output [31:0] Y;

	wire [31:0] S1,S2,S3,S4,S5;
	
	assign S1=(B[4]==1)?{A[15:0],16'd0}:A;
	assign S2=(B[3]==1)?{S1[23:0],8'd0}:S1;
	assign S3=(B[2]==1)?{S2[27:0],4'd0}:S2;
	assign S4=(B[1]==1)?{S3[29:0],2'd0}:S3;
	assign Y=(B[0]==1)?{S4[30:0],1'b0}:S4;

endmodule

module RSFT(Y,A,B);
	input  [31:0] A,B;
	output [31:0] Y;

	wire [31:0] S1,S2,S3,S4,S5;

	assign S1=(B[4]==1)?{16'd0,A[31:16]}:A;
	assign S2=(B[3]==1)? {8'd0,S1[31:8]}:S1;
	assign S3=(B[2]==1)? {4'd0,S2[31:4]}:S2;
	assign S4=(B[1]==1)? {2'd0,S3[31:2]}:S3;
	assign Y=(B[0]==1)? {1'b0,S4[31:1]}:S4;

endmodule

module ARSFT(Y,A,B);
	input  [31:0] A,B;
	output [31:0] Y;

	wire [31:0] S1,S2,S3,S4,S5;
	wire [15:0] S6;

	assign S6=(A[31]==1)?16'hFFFF:16'd0;//S6= xxxx xxxx xxxx xxxx  xxxx xxxx xxxx xxxx

	assign S1=(B[4]==1)?{S6,A[31:16]}:A;
	assign S2=(B[3]==1)?{S6[7:0],S1[31:8]}:S1;
	assign S3=(B[2]==1)?{S6[3:0],S2[31:4]}:S2;
	assign S4=(B[1]==1)?{S6[1:0],S3[31:2]}:S3;
	assign Y =(B[0]==1)?{S6[0],S4[31:1]}:S4;

endmodule

	/*always@(*)
	begin

		if(B[4]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^4=16 10000=16
			S1={S6,A[31:16]};		// xxxx xxxx xxxx xxxx  1111 1111 1111 1111   
		else
			S1=A;

		if(B[3]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^3=8 1000=8
			S2={S6[7:0],S1[31:8]};	// xxxx xxxx 1111 1111  1111 1111 1111 1111 
		else
			S2=S1;

		if(B[2]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^2=4 100=4
			S3={S6[3:0],S2[31:4]};	// xxxx 1111 1111 1111  1111 1111 1111 1111 
		else
			S3=S2;
		if(B[1]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^1=2 10=2
			S4={S6[1:0],S3[31:2]};  // xx11 1111 1111 1111  1111 1111 1111 1111 
		else
			S4=S3;
		if(B[0]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^0=1 1=1
			Y={S6[0],S4[31:1]};	// x111 1111 1111 1111  1111 1111 1111 1111 
		else
			Y=S4;
	end */
		/*always@(*)
	begin

		if(B[4]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^4=16 10000=16
			S1={16'd0,A[31:16]};		// 1111 1111 1111 1111  0000 0000 0000 0000 
		else
			S1=A;

		if(B[3]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^3=8 1000=8
			S2={8'd0,S1[31:8]};		// 1111 1111 1111 1111  1111 1111 0000 0000 
		else
			S2=S1;

		if(B[2]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^2=4 100=4
			S3={4'd0,S2[31:4]};		// 1111 1111 1111 1111  1111 1111 1111 0000 
		else
			S3=S2;
		if(B[1]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^1=2 10=2
			S4={2'd0,S3[31:2]};		// 1111 1111 1111 1111  1111 1111 1111 1100 
		else
			S4=S3;
		if(B[0]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^0=1 1=1
			S5={1'b0,S4[31:1]};		// 1111 1111 1111 1111  1111 1111 1111 1110 
		else
			S5=S4;
	end*/
		/*always@(*)
	begin

		if(B[4]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^4=16 10000=16
			S1={A[15:0],16'd0};		// 1111 1111 1111 1111  0000 0000 0000 0000 
		else
			S1=A;

		if(B[3]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^3=8 1000=8
			S2={S1[23:0],8'd0};		// 1111 1111 1111 1111  1111 1111 0000 0000 
		else
			S2=S1;

		if(B[2]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^2=4 100=4
			S3={S2[27:0],4'd0};		// 1111 1111 1111 1111  1111 1111 1111 0000 
		else
			S3=S2;
		if(B[1]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^1=2 10=2
			S4={S3[29:0],2'd0};		// 1111 1111 1111 1111  1111 1111 1111 1100 
		else
			S4=S3;
		if(B[0]==1)					// 1111 1111 1111 1111  1111 1111 1111 1111   2^0=1 1=1
			S5={S4[30:0],1'b0};		// 1111 1111 1111 1111  1111 1111 1111 1110 
		else
			S5=S4;
	end*/